* AD8138 SPICE Macro-model
* Description: Amplifier
* Generic Desc: Low distortion diff I/O amp - 500 MHz
* Developed by: JG/ADI, TRW/ADI
* Revision History: 08/10/2012 - Updated to new header style
* 5.0 (11/2002)
* Copyright 1999, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*     vnoise, not included in this version
*     inoise, not included in this version
*     distortion is not characterized
*     cmrr is not  characterized in this version.
*
* Parameters modeled include:
*     closed loop gain and phase vs bandwidth
*     output current and voltage limiting
*     offset voltage (is  non-static, will  vary with gain)
*     ibias (again, is static, will not vary with vcm)
*     slew rate and step response performance
*     (slew rate is based on 10-90% of step response)
*     current on output will be reflected to the supplies
*     Vocm is variable and include input typical offset
*
* END Notes:
*
* Node assignments
*                 non-inverting input
*                 | inverting input
*                 | | positive supply
*                 | | |  negative supply
*                 | | |  |  output positive
*                 | | |  |  |   output negative
*                 | | |  |  |   |   vocm input
*                 | | |  |  |   |   |
*.SUBCKT ad8138  3a 9 99 50 71b 71  110
.SUBCKT ad8138  +IN -IN VS+ VS- +OUT -OUT  VOCM
****************************input stage*******************************************


*****positive input left side*****

I1 VS+ 5 .4E-3
Q1 VS- 2 5 QX
vos +IN 2 -1.95E-3

**RAIL CLIPING****

Dlim+ 75 14b dx
Vlim+ VS+ 14b 2.1
Dlim 14c 75 dx
Vlim 14c  VS- 2.1
Dlim- 13b 76 DX
Vlim- 13b VS- 2.1
Dlim-B 76 13C dx
Vlim-B VS+ 13C 2.1

** VOCM INPUT RAIL CLIPING****

DOCMa 100 100A dx
VOCMa VS+ 100A 1.899
DOCMb 100b 100 DX
VOCMb 100b VS- 1.899

*****negative input right side*****

I2 VS+ 6 .4E-3
Q2 VS- -IN 6 QX

***********Input capacitance/impedance*******

Cin +IN -IN 1p

***************************************pole, zero pole stage********************************************

G1 13 14 5 6 5e-3
c1 14 13 1.7p
c2 13 98 .6p
c3 14 98 .6p
r11 13 98 250k
r12 14 98 250k

*********pole zero stage( POSITIVE SIDE)*******

gp1 0 75 14 98 1
RP1 75 0 1
CP1 75 0 .38E-9

*********pole zero stage( NEGATIVE SIDE)*******

gp2 0 76 13 98 1
RP2 76 0 1
CP2 76 0 .38E-9

**********output stage Negative side*************

D17 76 84 DX
VO1  84 70 .177V
VO2  70 85 .177V
D16 85 76  DX
G30 70 99c VS+ 76  91E-3
G31 98c 70 76 VS-  91E-3
RO30 70 99c 11
RO31 98c 70 11
VIOUT1 VS+ 99c 0V
VIOUT2 VS- 98c 0V
VIOUT3 70 -OUT 0V

********** Output Stage Positive side *************

D17b 75 84b DX
VO1b  84b 70b .177V
VO2b  70b 85b .177V
D16b 85b 75  DX
G30b 70b 99d VS+ 75  91E-3
G31b 98d 70b 75 VS-  91E-3
RO30b 70b 99d 11
RO31b 98d 70b 11
VIOUTB1 VS+ 99d 0V
VIOUTB2 98d VS- 0V
VIOUTB3 70b +OUT 0V

*********VOCM STAGE*************************

Gocm_a 0 75 VOCM 0 1
Gocm_b 0 76 VOCM 0 1
Rocm1 VS+ 100 400k
Rocm2 100 VS- 400k
Voffset 100 VOCM -1E-3

********CURRENT MIRROR TO SUPPLIES POSITVIE SIDE*********

FO1 0 VS+ poly(2) VIOUT1 VI1 -19.803E-3 1 -1
FO2 0 VS- poly(2) VIOUT2 VI2 -19.803E-3 1 -1
FO3 0 400 VIOUT1 1
VI1 401 0 0
VI2 0 402 0
DM1 400 401 DX
DM2 402 400 DX

********CURRENT MIRROR TO SUPPLIES NEGATIVE SIDE*********

FO1B 0 VS+ poly(2) VIOUTB1 VIB1 -19.803E-3 1 -1
FO2B 0 VS- poly(2) VIOUTB2 VIB2 -19.803E-3 1 -1
FO3B 0 400B VIOUTB1 1
VIB1 401B 0 0
VIB2 0 402B 0
DMB1 400B 401B DX
DMB2 402B 400B DX

***  Reference Stage

Eref 98 0 poly(2) VS+ 0 VS- 0 0 0.5 0.5



.MODEL QX PNP (BF=228.57 Is=1E-15)
.MODEL DX D(IS=1E-15)
.ENDS






